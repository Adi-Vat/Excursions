package instruction_set;
	typedef enum logi[7:0]
	{
		NOP, // NO OPERATION
		LDD, // LOAD DIRECLTY INTO REGISTER <REG> FROM <MEMORY/REG>
		LDD_I, // LOAD DIRECTLY INTO REGISTER <REG> FROM >VALUE>
		LDR, // LOAD INTO REGISTER <REG> DATA AT MEMORY LOCATION IN <MEMORY/REG>
		STR, // STORE INTO <MEMORY> DATA FROM <REG>
		STR_I, // STORE
		ADC, // ADD WITH CARRY ACC AND <REG/VALUE> STORE INTO ACC
		ADC_I,
		SUB, // SUBTRACT ACC AND <REG/VALUE> STORE INTO ACC
		SUB_I,
		INC, // INCREMENT <REG>
		DEC, // DECREMENT <REG>
		ROL, // ROTATE LEFT <REG>
		ROR, // ROTATE RIGHT <REG>
		SLL, // SHIFT LEFT LOGICAL <REG>
		SLA, // SHIFT LEFT ARITHMETIC <REG>
		SRL, // SHIFT RIGHT LOGICAL <REG>
		SRA, // SHIFT RIGHT ARITHMETIC <REG>
		PSH, // PUSH <REG> TO STACK
		POP, // POP STACK ONTO <REG>
		JMP, // JUMP TO <VAL>
		CMP, // COMPARE <REG> WITH ACC
		CMP_I,
		JZ, // JUMP TO <VAL> IF ZERO FLAG IS SET
		JNZ, // JUMP TO <VAL> IF ZERO FLAG IS NOT SET
		JN, // JUMP TO <VAL> IF NEGATIVE FLAG IS SET
		SB, // SET AT <MEMORY/REG> BIT NUMBER <VAL> TO 1
		CB // CLEAR AT <MEMORY/REG> BIT NUMBER <VAL> TO 0
	} OPCODES;
endpackage